module dataPath() ;
	


endmodule
