//James Jhong
//Jean Kim
//EE469 Lab 2
//1/18/2022

//This module is a 1 bit slice of the alu, a 4:1 mux.
//It can handle 4 operations, addition, subtraction, AND and OR.
//It has two inputs A and B. 

module alu_1bit_slice(a, b, cin, co, control, out);
	//add or subtract, Cin, Cout, uses the 2 x 1 mux to determine which one
		
endmodule
